module UART_Tx
(
    input logic clk, reset,
    input logic transmit,
    input logic [31:0] tx_bits,
    output logic output_stream
);

endmodule: UART_Tx
