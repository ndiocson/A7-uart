module UART_Rx 
(   
    input logic clk, reset,
    input logic input_stream,
    output logic [31:0] rx_bits
);

endmodule: UART_Rx
